`include "tmod_master.sv"
`include "tmod_slave.sv"
`include "temp_sensor.sv"
