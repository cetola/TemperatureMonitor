`include "tmod-master.sv"
`include "tmod-slave.sv"
`include "temp-sensor.sv"