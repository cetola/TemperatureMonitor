`include "defs.sv"
module temp_sensor(input logic clk, input logic reset, output logic tick, output logic[7:0] temp);
    
endmodule